module inv_kicad_sch(
    output Y,
    input A);

    NOT U4(A, Y);
endmodule
