module inv_kicad_sch(
    input A,
    output Y);

    // TBD wires

    74LS04 U4(/* */);
endmodule
