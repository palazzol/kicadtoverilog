module inv(
    output Y,
    input A);

    NOT U3(.A(A), .Y(Y));
endmodule
