module inv_kicad_sch(
    output Y,
    input A);

    NOT U3(A, Y);
endmodule
