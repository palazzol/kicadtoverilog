module inv_kicad_sch(
    output Y,
    input A);

    wire w1;
    wire w2;

    NOT U4(/* */);
endmodule
